module processor(
    input wire clk,
    input wire rst
);
endmodule

module alu(

);
endmodule

module load(

);
endmodule

module store(

);
endmodule